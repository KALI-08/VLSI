class transactions;
  rand bit clk,reset;
  bit [7:0]out;
endclass
