module top_module (
    output reg out);
assign out=1'b0;
endmodule
