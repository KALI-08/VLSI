interface alu_if(input logic clk);
  logic [3:0] a, b;
    logic [1:0] op;
  logic [3:0] result;

endinterface
