interface operation;
  logic a,b;
  logic sum,carry;
endinterface
