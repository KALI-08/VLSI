interface intf;
  logic clk,reset,w_en,r_en;
  logic [7:0]data_in;
  logic [7:0]data_out;
  logic full,empty;
endinterface
  
