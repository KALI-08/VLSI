interface dff_intf(input logic clk);
  logic rst;
  logic d;
  logic q;
endinterface
