interface operation;
  logic clk,reset;
  logic [7:0]out;
endinterface
