// Code your design here
module or_gate(
  input a,b,
  output c);
  or(c,a,b);
endmodule
