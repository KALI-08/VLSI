module xnor_gate(
  input x,y,
  output z);
  xnor (z,x,y);
endmodule
