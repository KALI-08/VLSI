// Code your design here
module nor_gate(
  input a,b,
  output c);
  nor (c,a,b);
endmodule
