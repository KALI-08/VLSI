// Code your design here
module and_gate(
  input A,B,
  output Y);
  and(Y,A,B);
endmodule
