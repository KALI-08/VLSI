// Code your design here
module xor_gate(
  input a,b,
  output c);
  xor (c,a,b);
endmodule
